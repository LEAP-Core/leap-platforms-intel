//
// Copyright (c) 2016, Intel Corporation
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
//
// Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation
// and/or other materials provided with the distribution.
//
// Neither the name of the Intel Corporation nor the names of its contributors
// may be used to endorse or promote products derived from this software
// without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF
// SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS
// INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN
// CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.

`include "cci_mpf_if.vh"
`include "cci_mpf_shim_edge.vh"

//
// This is a mandatory connection at the head of an MPF pipeline.
// It canonicalizes input and output and manages the flow of data through
// MPF.
//

module cci_mpf_shim_edge_afu
  #(
    parameter N_WRITE_HEAP_ENTRIES = 0,

    // Enforce write/write and write/read ordering with cache lines?
    parameter ENFORCE_WR_ORDER = 0
    )
   (
    input  logic clk,

    // Connection toward the FIU (the end of the MPF pipeline nearest the AFU)
    cci_mpf_if.to_fiu fiu,

    // External connections to the AFU
    cci_mpf_if.to_afu afu,

    // Interface to the MPF FIU edge module
    cci_mpf_shim_edge_if.edge_afu fiu_edge
    );

    logic reset;
    assign reset = fiu.reset;

    // Have the AFU come out of reset a cycle late both to allow the MPF
    // distributed reset tree to complete and to put the AFU in a separate
    // reset domain.
    initial
    begin
        afu.reset = 1'b1;
    end

    always @(posedge clk)
    begin
        afu.reset <= fiu.reset;
    end


    //
    // Save write data as it arrives from the AFU in a heap here.  Use
    // the saved values as requests exit MPF toward the FIU.  This has
    // multiple advantages:
    //
    //   - Internal buffer space inside MPF pipelines is greatly reduced
    //     since the wide request channel 1 data bus is eliminated.
    //
    //   - Multi-beat write requests are easier to handle.  The code
    //     here will send only one write request through MPF.  The remaining
    //     beats are saved in the heap here and regenerated when the
    //     control packet exits MPF.
    //
    typedef logic [$clog2(N_WRITE_HEAP_ENTRIES)-1 : 0] t_write_heap_idx;

    logic wr_heap_alloc;
    logic wr_heap_not_full;
    t_write_heap_idx wr_heap_enq_idx;
    t_cci_clNum wr_heap_enq_clNum;

    cci_mpf_prim_heap_ctrl
      #(
        .N_ENTRIES(N_WRITE_HEAP_ENTRIES),
        // Leave space both for the almost full threshold and a full
        // multi-line packet.  To avoid deadlocks we never signal a
        // transition to almost full in the middle of a packet so must
        // be prepared to absorb all flits.
        .MIN_FREE_SLOTS(CCI_TX_ALMOST_FULL_THRESHOLD +
                        CCI_MAX_MULTI_LINE_BEATS + 1)
        )
      wr_heap_ctrl
       (
        .clk,
        .reset,

        // Add entries to the heap as writes arrive from the AFU
        .enq(wr_heap_alloc),
        .notFull(wr_heap_not_full),
        .allocIdx(wr_heap_enq_idx),

        // Free entries as writes leave toward the FIU.
        .free(fiu_edge.free),
        .freeIdx(fiu_edge.freeidx)
        );


    //
    // The heap holding write data is in the FIU edge module.
    //
    assign fiu_edge.wen = cci_mpf_c1TxIsWriteReq(afu.c1Tx);
    assign fiu_edge.widx = wr_heap_enq_idx;
    assign fiu_edge.wclnum = wr_heap_enq_clNum;
    assign fiu_edge.wdata = afu.c1Tx.data;


    // ====================================================================
    //
    //   AFU edge flow
    //
    // ====================================================================

    logic afu_wr_packet_active;
    logic afu_wr_sticky_full;
    logic afu_wr_eop;

    assign wr_heap_alloc = cci_mpf_c1TxIsWriteReq(afu.c1Tx) && afu_wr_eop;

    logic afu_wr_almost_full;
    assign afu_wr_almost_full = fiu.c1TxAlmFull || ! wr_heap_not_full;

    // All but write requests flow straight through. The c1Tx channel needs
    // to be registered in this module due to the logic that drops all but
    // one flit from a multi-beat write.  If read/write order is being
    // enforced than add the same register latency for c0Tx.
    generate
        if (ENFORCE_WR_ORDER)
        begin : wr_order
            always_ff @(posedge clk)
            begin
                fiu.c0Tx <= cci_mpf_updC0TxCanonical(afu.c0Tx);
            end
        end
        else
        begin : no_wr_order
            assign fiu.c0Tx = cci_mpf_updC0TxCanonical(afu.c0Tx);
        end
    endgenerate

    assign fiu.c2Tx = afu.c2Tx;

    //
    // Register almost full signals before they reach the AFU.  MPF modules
    // must accommodate the extra cycle of buffering that may be needed
    // as a result of signalling almost full a cycle late.
    //
    always_ff @(posedge clk)
    begin
        if (reset)
        begin
            afu.c0TxAlmFull <= 1'b1;
            afu.c1TxAlmFull <= 1'b1;
            afu_wr_sticky_full <= 1'b0;
        end
        else
        begin
            afu.c0TxAlmFull <= fiu.c0TxAlmFull;

            // Never signal almost full in the middle of a packet. Deadlocks
            // can result since the control flit is already flowing through MPF.
            afu.c1TxAlmFull <= afu_wr_almost_full &&
                                   (! afu_wr_packet_active || afu_wr_sticky_full);

            // afu_wr_sticky_full goes high as soon as afu_wr_almost_full is
            // asserted and no packet is in flight.  It stays high until
            // afu_wr_almost_full is no longer asserted.
            if (! afu_wr_almost_full)
            begin
                afu_wr_sticky_full <= 1'b0;
            end
            else if (afu_wr_almost_full && ! afu_wr_packet_active)
            begin
                afu_wr_sticky_full <= 1'b1;
            end
        end
    end

    assign afu.c0Rx = fiu.c0Rx;
    assign afu.c1Rx = fiu.c1Rx;

    //
    // The CCI spec. allows both address and cl_len of non-sop flits in a
    // multi-beat packet to be don't care, which is rather annoying.
    // Register the sop values and add a mux to recover them.
    //
    t_cci_clLen c1tx_sop_clLen;
    t_cci_clAddr c1tx_sop_clAddr;

    always_ff @(posedge clk)
    begin
        if (afu.c1Tx.hdr.base.sop == 1'b1)
        begin
            c1tx_sop_clLen <= afu.c1Tx.hdr.base.cl_len;
            c1tx_sop_clAddr <= afu.c1Tx.hdr.base.address;
        end
    end

    // Generate canonical c1Tx, including cl_len and address.
    t_if_cci_mpf_c1_Tx afu_canon_c1Tx;

    always_comb
    begin
        afu_canon_c1Tx = cci_mpf_updC1TxCanonical(afu.c1Tx);

        if (! afu.c1Tx.hdr.base.sop)
        begin
            afu_canon_c1Tx.hdr.base.cl_len = c1tx_sop_clLen;
            afu_canon_c1Tx.hdr.base.address = c1tx_sop_clAddr;
        end
    end


    always_ff @(posedge clk)
    begin
        fiu.c1Tx <= cci_mpf_updC1TxCanonical(afu_canon_c1Tx);

        // The cache line's value stored in fiu.c1Tx.data is no longer needed
        // in the pipeline.  Store 'x but use the low bits to hold the
        // local heap index.
        fiu.c1Tx.data <= 'x;
        fiu.c1Tx.data[$clog2(N_WRITE_HEAP_ENTRIES) - 1 : 0] <= wr_heap_enq_idx;

        // Multi-beat write request?  Only the start of packet beat goes
        // through MPF.  The rest are buffered in wr_heap here and the
        // packets will be regenerated when the sop packet exits.
        //
        // Only pass requests that are either the end of a write or
        // that aren't writes.
        if (cci_mpf_c1TxIsWriteReq_noCheckValid(afu_canon_c1Tx))
        begin
            // Wait for the final flit to arrive and be buffered, thus
            // guaranteeing that all the data is ready to be written
            // as the packet exits to the FIU.
            fiu.c1Tx.valid <= afu_canon_c1Tx.valid &&
                              (wr_heap_enq_clNum == afu_canon_c1Tx.hdr.base.cl_len);

            fiu.c1Tx.hdr.base.sop <= 1'b1;
        end
    end


    //
    // Validate request.  All the remaining code is just validation that
    // multi-beat requests are formatted properly.
    //

    cci_mpf_prim_track_multi_write
      afu_wr_track
       (
        .clk,
        .reset,
        .c1Tx(afu_canon_c1Tx),
        .c1Tx_en(1'b1),
        .eop(afu_wr_eop),
        .packetActive(afu_wr_packet_active),
        .nextBeatNum(wr_heap_enq_clNum)
        );

    t_cci_clLen afu_wr_prev_cl_len;

    always_ff @(posedge clk)
    begin
        if (reset)
        begin
            // Nothing
        end
        else
        begin
            if (cci_mpf_c0TxIsReadReq(afu.c0Tx))
            begin
                assert((afu.c0Tx.hdr.base.address[1:0] & afu.c0Tx.hdr.base.cl_len) == 2'b0) else
                    $fatal("cci_mpf_shim_edge_connect: Multi-beat read address must be naturally aligned");
            end

            if (cci_mpf_c1TxIsWriteReq(afu_canon_c1Tx))
            begin
                assert(afu.c1Tx.hdr.base.sop != afu_wr_packet_active) else
                    if (! afu.c1Tx.hdr.base.sop)
                        $fatal("cci_mpf_shim_edge_connect: Expected SOP flag on write");
                    else
                        $fatal("cci_mpf_shim_edge_connect: Wrong number of multi-beat writes");

                if (afu.c1Tx.hdr.base.sop)
                begin
                    assert ((afu.c1Tx.hdr.base.address[1:0] & afu_canon_c1Tx.hdr.base.cl_len) == 2'b0) else
                        $fatal("cci_mpf_shim_edge_connect: Multi-beat write address must be naturally aligned");
                end
                else
                begin
                    assert (afu_wr_prev_cl_len == afu_canon_c1Tx.hdr.base.cl_len) else
                        $fatal("cci_mpf_shim_edge_connect: cl_len must be the same in all beats of a multi-line write");
                end

                afu_wr_prev_cl_len <= afu_canon_c1Tx.hdr.base.cl_len;
            end
        end
    end

endmodule // cci_mpf_shim_edge_afu

