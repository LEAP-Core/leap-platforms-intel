//
// MPF's view of CCI expressed as a SystemVerilog interface.
//

`ifndef CCI_MPF_IF_VH
`define CCI_MPF_IF_VH

import cci_mpf_if_pkg::*;

`ifdef USE_PLATFORM_CCI_S
import ccis_if_pkg::*;
`endif

`ifdef USE_PLATFORM_CCI_P
import ccip_if_pkg::*;
`endif

// Global log file handle
int cci_mpf_if_log_fd = -1;

interface cci_mpf_if
  #(
    parameter ENABLE_LOG = 0,        // Log events for this instance?
    parameter LOG_NAME = "cci_mpf_if.tsv"
    )
   (
    input logic clk
    );

    // Reset flows from QLP to AFU
    logic              reset_n;

    // Requests to QLP.  All objects are outputs flowing toward QLP except
    // the almost full ports, which provide flow control.
    t_if_cci_mpf_c0_Tx c0Tx;
    logic              c0TxAlmFull;

    t_if_cci_mpf_c1_Tx c1Tx;
    logic              c1TxAlmFull;

    // Responses from QLP.  All objects are inputs from the QLP and flow
    // toward the AFU.  There is no flow control.  The AFU must be prepared
    // to receive responses for all in-flight requests.
    t_if_cci_c0_Rx     c0Rx;
    t_if_cci_c1_Rx     c1Rx;

    // Port directions for connections in the direction of the QLP (platform)
    modport to_qlp
      (
       input  reset_n,

       output c0Tx,
       input  c0TxAlmFull,

       output c1Tx,
       input  c1TxAlmFull,

       input  c0Rx,
       input  c1Rx
       );

    // Port directions for connections in the direction of the AFU (user code)
    modport to_afu
      (
       output reset_n,

       input  c0Tx,
       output c0TxAlmFull,

       input  c1Tx,
       output c1TxAlmFull,

       output c0Rx,
       output c1Rx
       );


    // ====================================================================
    //
    // Snoop equivalents of the above interfaces: all the inputs and none
    // of the outputs.
    //
    // ====================================================================

    modport to_qlp_snoop
      (
       input  reset_n,

       input  c0TxAlmFull,
       input  c1TxAlmFull,

       input  c0Rx,
       input  c1Rx
       );

    modport to_afu_snoop
      (
       input  reset_n,

       input  c0Tx,
       input  c1Tx
       );


    // ====================================================================
    //
    //   Debugging
    //
    // ====================================================================

`ifdef CCI_SIMULATION

`include "cci_mpf_if_dbg.vh"

`endif

endinterface

`endif //  CCI_MPF_IF_VH
